netcdf foo {  // an example netCDF specification in CDL

              types:
                  ubyte enum enum_t {Clear = 0, Cumulonimbus = 1, Stratus = 2};
                  opaque(11) opaque_t;
                  int(*) vlen_t;

              dimensions:
                   lat = 10, lon = 5, time = unlimited ;
                   height = 100 ;

              variables:
                   ubyte   tag;
                   double  p(time,lat,lon);
                   long    rh(time,lat,lon);
                   string  country(time,lat,lon);
                   long    lat(lat), lon(lon), time(time);
                   float   Z(time,lat,lon), t(time,lat,lon);


                   // variable attributes
                   :untyped_global_attribute = "global";
                   lat:long_name = "latitude";
                   lat:units = "degrees_north";
                   lon:long_name = "longitude";
                   lon:units = "degrees_east";
                   time:units = "seconds since 1992-1-1 00:00:00";

                   // typed variable attributes
                   string Z:units = "geopotential meters";
                   float Z:valid_range = 0., 5000.;
                   double p:_FillValue = -9999.;
                   long rh:_FillValue = -1;
                   vlen_t :globalatt = {17, 18, 19};
              data:
                   lat   = 0, 10, 20, 30, 40, 50, 60, 70, 80, 90;
                   lon   = -140, -118, -96, -84, -52;
              group: g {
              types:
                  compound cmpd_t { vlen_t f1; enum_t f2;};
              } // group g
              group: h {
              variables:
                   /g/cmpd_t  compoundvar;
             data:
	              compoundvar = { {3,4,5}, enum_t.Stratus } ;
    } // group h
}
